library verilog;
use verilog.vl_types.all;
entity Adder16_TB is
end Adder16_TB;
